##INPUTS
set_property PACKAGE_PIN K18 [get_ports {UP}]
set_property IOSTANDARD LVCMOS33 [get_ports {UP}]

set_property PACKAGE_PIN P16 [get_ports {DOWN}]
set_property IOSTANDARD LVCMOS33 [get_ports {DOWN}]

set_property PACKAGE_PIN K19 [get_ports {RESET}]
set_property IOSTANDARD LVCMOS33 [get_ports {RESET}]

set_property PACKAGE_PIN L16 [get_ports {CLOCK}]
set_property IOSTANDARD LVCMOS33 [get_ports {CLOCK}]

##LEDS
set_property PACKAGE_PIN M14 [get_ports {LEDS[0]}]
set_property IOSTANDARD LVCMOS33 [get_ports {LEDS[0]}]

set_property PACKAGE_PIN M15 [get_ports {LEDS[1]}]
set_property IOSTANDARD LVCMOS33 [get_ports {LEDS[1]}]

set_property PACKAGE_PIN G14 [get_ports {LEDS[2]}]
set_property IOSTANDARD LVCMOS33 [get_ports {LEDS[2]}]

set_property PACKAGE_PIN D18 [get_ports {LEDS[3]}]
set_property IOSTANDARD LVCMOS33 [get_ports {LEDS[3]}]